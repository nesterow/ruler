module main

import rest

fn main() {
	rest.serve()!
}
