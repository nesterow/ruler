module task

fn test_task_service() {}
