module task

pub struct TaskService {}
