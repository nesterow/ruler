module dto

pub struct UpdateTaskIndexDTO {
pub:
	worker_name string
}
